interface LeadingZeroCounter;
	method Bool read_rs1();
	method Action load_rs1(Bit#(8) newval);
	method Bit#(8) read_count();
	method Action increment_count();
	method Bit#(8) read_rs1value();
	method Action leftshift_rs1(Bit#(8) shiftvalue);
endinterface

(*synthesize*)
module mkLeadingZeroCounter(LeadingZeroCounter);
	Reg#(Bit#(8)) rg_rs1 <- mkRegU();
	Reg#(Bit#(8)) count <- mkReg(0);
	method Action load_rs1(Bit#(8) newval);
		rg_rs1 <= newval;
	endmethod
	method Bit#(8) read_rs1value();
		return rg_rs1;
	endmethod
	method Bool read_rs1();
		if(rg_rs1[7]==1) return True;
		else return False;
	endmethod
	method Bit#(8) read_count();
		return count;
	endmethod
	method Action increment_count();
		count <= count + 1;
	endmethod
	method Action leftshift_rs1(Bit#(8) shiftvalue);
		rg_rs1 <= rg_rs1 << shiftvalue;
	endmethod
endmodule
